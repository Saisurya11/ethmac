typedef uvm_sequencer#(eth_frame) phy_rx_sqr;